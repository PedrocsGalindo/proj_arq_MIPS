module PCAdder (
    input wire [31:0] pc_in,   // Entrada: valor atual do PC
    output wire [31:0] pc_out  // Saída: PC atualizado
);
    assign pc_out = pc_in + 4; // Incrementa o PC em 4
endmodule
